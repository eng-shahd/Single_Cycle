library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

   --> funct codes <--
--------------------------------
-- add         		  | 100000 |
-- subtract    		  | 100010 |
-- and         		  | 100100 |
-- or          		  | 100101 |
-- nor         		  | 100111 |
-- shift_left  		  | 000000 |
-- shift_right 		  | 000010 |
-- set_is_less_than   | 101010 |
--------------------------------

entity ALUControl is
  port(
    ALUOp      : in  std_logic_vector(1 downto 0);
    funct      : in  std_logic_vector(5 downto 0);
    ALUControl : out std_logic_vector(3 downto 0) );
end entity;

architecture Behavior of ALUControl is
begin

  process(ALUOp, funct)
  begin
    case ALUOp is

      -- LW, SW => ADD 
      when "00" =>
        ALUControl <= "0000";

      -- BEQ => SUB
      when "01" =>
        ALUControl <= "0001";

      -- R-type
      when "10" =>
        case funct is
          when "100000" => ALUControl <= "0000"; -- add
          when "100010" => ALUControl <= "0001"; -- sub
          when "100100" => ALUControl <= "0010"; -- and
          when "100101" => ALUControl <= "0011"; -- or
          when "100111" => ALUControl <= "0100"; -- nor
          when "000000" => ALUControl <= "0101"; -- sll
          when "000010" => ALUControl <= "0110"; -- srl
	  when "101010" => ALUControl <= "0111"; -- slt
          when others   => ALUControl <= "1111"; -- undefined
        end case;

      when others =>
        ALUControl <= "1111";

    end case;
  end process;

end architecture;
